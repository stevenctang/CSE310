module main();// Always have to call your module something
	initial	  
	begin
	$display("Steven");
	end
endmodule// Always have to have the end module, everything goes inside of here
